../Aufgabe02/aluCtrlExt.vhd