../../../Blatt05/praxis/Aufgabe03/proc_config.vhd