../../../Blatt09/praxis/Aufgabe02/proc_config.vhd