../../../Blatt03/praxis/Aufgabe03/bin2Char.vhd