../../../Blatt07/praxis/Aufgabe02/alu_1bit.vhd