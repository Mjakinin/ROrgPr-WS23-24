../../../Blatt08/praxis/Aufgabe02/mipsISA.vhd