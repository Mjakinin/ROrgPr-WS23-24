../../../Blatt08/praxis/Aufgabe02/alu_1bit.vhd