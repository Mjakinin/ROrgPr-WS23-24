../../../Blatt07/praxis/Aufgabe02/adder_1bit.vhd