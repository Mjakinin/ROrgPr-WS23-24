../../../Blatt09/praxis/Aufgabe02/mipsCtrlFsm.vhd