../Aufgabe02/alu_1bit.vhd