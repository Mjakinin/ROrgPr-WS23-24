../../../Blatt06/praxis/Aufgabe02/addrDecoder.vhd