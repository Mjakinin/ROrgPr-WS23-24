../../../Blatt07/praxis/Aufgabe03/mipsAlu.vhd