../Aufgabe02/addrDecoder.vhd