../../../Blatt04/praxis/Aufgabe01/signExtend.vhd