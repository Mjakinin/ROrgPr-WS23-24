../../../Blatt04/praxis/Aufgabe02/leftShifter.vhd