../../../Blatt08/praxis/Aufgabe01/mipsISA.vhd