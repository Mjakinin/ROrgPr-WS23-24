../../../Blatt06/praxis/Aufgabe03/regFile.vhd