../../../Blatt00/praxis/Aufgabe01/or2.vhd