../../../Blatt01/praxis/Aufgabe01/xor2.vhd