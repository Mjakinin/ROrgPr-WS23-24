../../../Blatt07/praxis/Aufgabe01/aluCtrl.vhd