library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;

library std;
use std.textio.all;

library work;
use work.mipsISA.all;


entity aluCtrlExt_tb is
end aluCtrlExt_tb;

architecture behavioral of aluCtrlExt_tb is

begin

    -- Beschreibung der Testbench ergänzen

    -- Ihr könnt ein `report "CI: All good." severity note;` einfügen (nur im Erfolgsfall),
    -- damit die automatischen Tests auch mit eurer Testbench funktionieren.
end behavioral;
