../../../Blatt05/praxis/Aufgabe02.2/reg.vhd