../Aufgabe01/mipsISA.vhd