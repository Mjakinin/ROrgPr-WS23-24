../../praxis/Aufgabe01/mipsCtrl.vhd