../Aufgabe02/adder_1bit.vhd